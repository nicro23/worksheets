
module adder(input a,input b, input cin, output s, output cout)


endmodule

module multi_adder(input a0, input a1,input a2, input a3, input b0, input b1, input b2, input b3, input cin,output s0, output s1, output s2, output s3, output cout)

begin
    
end
endmodule